// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

interface synapse_if
( input clk
, input reset
);
  // --------------------------------------------------------------------
  int weight = 3;
  wire spike;

// --------------------------------------------------------------------
endinterface
