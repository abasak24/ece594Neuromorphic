// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

interface synapse_if
( input clk
, input reset
);
  // --------------------------------------------------------------------
  int weight = 1;
  wire spike;

// --------------------------------------------------------------------
endinterface
