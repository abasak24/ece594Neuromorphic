localparam neuron_config_t CFG = '{1, 0, 0, 1, ALPHA};

localparam int S[T][N] = 
'{ '{18, 20, 23, 19, 20, 21, 16, 18, 19, 15, 23, 17, 18, 18, 22, 19, 18, 19, 22, 22, 25, 23, 22, 17, 20, 25, 18, 15, 23, 18, 19, 20}};

defparam block[0].nb.neuron[0].syn.SPIKE = {{0, 1}, {0, 2}, {0, 3}, {0, 5}, {0, 6}, {0, 8}, {0, 11}, {0, 12}, {0, 13}, {0, 14}, {0, 15}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 23}, {0, 24}};
defparam block[0].nb.neuron[1].syn.SPIKE = {{0, 0}, {0, 3}, {0, 4}, {0, 5}, {0, 7}, {0, 8}, {0, 12}, {0, 13}, {0, 15}, {0, 16}, {0, 18}, {0, 20}, {0, 21}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 26}, {0, 29}, {0, 31}};
defparam block[0].nb.neuron[2].syn.SPIKE = {{0, 0}, {0, 3}, {0, 8}, {0, 9}, {0, 10}, {0, 11}, {0, 12}, {0, 13}, {0, 14}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 27}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[3].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 5}, {0, 7}, {0, 9}, {0, 11}, {0, 13}, {0, 15}, {0, 16}, {0, 19}, {0, 20}, {0, 25}, {0, 26}, {0, 27}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[4].syn.SPIKE = {{0, 1}, {0, 3}, {0, 6}, {0, 8}, {0, 10}, {0, 12}, {0, 13}, {0, 14}, {0, 15}, {0, 17}, {0, 18}, {0, 20}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}, {0, 31}};
defparam block[0].nb.neuron[5].syn.SPIKE = {{0, 0}, {0, 1}, {0, 3}, {0, 6}, {0, 7}, {0, 8}, {0, 9}, {0, 10}, {0, 13}, {0, 14}, {0, 15}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 25}, {0, 26}, {0, 27}, {0, 30}};
defparam block[0].nb.neuron[6].syn.SPIKE = {{0, 0}, {0, 4}, {0, 5}, {0, 11}, {0, 12}, {0, 15}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 25}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[7].syn.SPIKE = {{0, 1}, {0, 3}, {0, 5}, {0, 9}, {0, 10}, {0, 11}, {0, 12}, {0, 14}, {0, 16}, {0, 18}, {0, 20}, {0, 21}, {0, 22}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}};
defparam block[0].nb.neuron[8].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 5}, {0, 10}, {0, 11}, {0, 13}, {0, 14}, {0, 15}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 31}};
defparam block[0].nb.neuron[9].syn.SPIKE = {{0, 2}, {0, 3}, {0, 5}, {0, 7}, {0, 10}, {0, 14}, {0, 15}, {0, 21}, {0, 22}, {0, 23}, {0, 25}, {0, 26}, {0, 28}, {0, 29}, {0, 31}};
defparam block[0].nb.neuron[10].syn.SPIKE = {{0, 2}, {0, 4}, {0, 5}, {0, 7}, {0, 8}, {0, 9}, {0, 11}, {0, 12}, {0, 14}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 21}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[11].syn.SPIKE = {{0, 0}, {0, 2}, {0, 3}, {0, 6}, {0, 7}, {0, 8}, {0, 10}, {0, 14}, {0, 16}, {0, 19}, {0, 20}, {0, 21}, {0, 24}, {0, 25}, {0, 26}, {0, 27}, {0, 29}};
defparam block[0].nb.neuron[12].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 6}, {0, 7}, {0, 10}, {0, 13}, {0, 14}, {0, 17}, {0, 20}, {0, 21}, {0, 22}, {0, 24}, {0, 27}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[13].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 3}, {0, 4}, {0, 5}, {0, 8}, {0, 12}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}};
defparam block[0].nb.neuron[14].syn.SPIKE = {{0, 0}, {0, 2}, {0, 4}, {0, 5}, {0, 7}, {0, 8}, {0, 9}, {0, 10}, {0, 11}, {0, 12}, {0, 15}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 25}, {0, 26}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[15].syn.SPIKE = {{0, 0}, {0, 1}, {0, 3}, {0, 4}, {0, 5}, {0, 6}, {0, 8}, {0, 9}, {0, 14}, {0, 16}, {0, 17}, {0, 19}, {0, 21}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[16].syn.SPIKE = {{0, 1}, {0, 2}, {0, 3}, {0, 7}, {0, 8}, {0, 10}, {0, 11}, {0, 15}, {0, 17}, {0, 19}, {0, 20}, {0, 22}, {0, 23}, {0, 25}, {0, 27}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[17].syn.SPIKE = {{0, 0}, {0, 2}, {0, 4}, {0, 5}, {0, 6}, {0, 8}, {0, 10}, {0, 12}, {0, 14}, {0, 15}, {0, 16}, {0, 18}, {0, 20}, {0, 21}, {0, 23}, {0, 24}, {0, 27}, {0, 28}, {0, 31}};
defparam block[0].nb.neuron[18].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 5}, {0, 6}, {0, 7}, {0, 8}, {0, 10}, {0, 13}, {0, 14}, {0, 17}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 23}, {0, 25}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[19].syn.SPIKE = {{0, 0}, {0, 2}, {0, 3}, {0, 5}, {0, 6}, {0, 8}, {0, 10}, {0, 11}, {0, 13}, {0, 14}, {0, 15}, {0, 16}, {0, 18}, {0, 20}, {0, 21}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[20].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 3}, {0, 4}, {0, 5}, {0, 6}, {0, 7}, {0, 11}, {0, 12}, {0, 13}, {0, 14}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 21}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 27}, {0, 28}, {0, 29}, {0, 30}};
defparam block[0].nb.neuron[21].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 5}, {0, 6}, {0, 7}, {0, 9}, {0, 10}, {0, 11}, {0, 12}, {0, 13}, {0, 14}, {0, 15}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 22}, {0, 23}, {0, 24}, {0, 27}, {0, 28}, {0, 29}};
defparam block[0].nb.neuron[22].syn.SPIKE = {{0, 1}, {0, 2}, {0, 4}, {0, 5}, {0, 6}, {0, 7}, {0, 8}, {0, 9}, {0, 10}, {0, 12}, {0, 13}, {0, 16}, {0, 18}, {0, 20}, {0, 21}, {0, 23}, {0, 24}, {0, 25}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[23].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 8}, {0, 9}, {0, 10}, {0, 16}, {0, 17}, {0, 18}, {0, 20}, {0, 21}, {0, 22}, {0, 26}, {0, 27}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[24].syn.SPIKE = {{0, 0}, {0, 1}, {0, 2}, {0, 4}, {0, 7}, {0, 8}, {0, 10}, {0, 11}, {0, 12}, {0, 13}, {0, 15}, {0, 17}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 26}, {0, 27}, {0, 28}, {0, 30}};
defparam block[0].nb.neuron[25].syn.SPIKE = {{0, 1}, {0, 2}, {0, 3}, {0, 4}, {0, 5}, {0, 6}, {0, 7}, {0, 8}, {0, 9}, {0, 10}, {0, 11}, {0, 13}, {0, 14}, {0, 15}, {0, 16}, {0, 18}, {0, 19}, {0, 20}, {0, 22}, {0, 26}, {0, 27}, {0, 28}, {0, 29}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[26].syn.SPIKE = {{0, 1}, {0, 3}, {0, 4}, {0, 5}, {0, 7}, {0, 9}, {0, 10}, {0, 11}, {0, 13}, {0, 14}, {0, 15}, {0, 19}, {0, 23}, {0, 24}, {0, 25}, {0, 27}, {0, 28}, {0, 30}};
defparam block[0].nb.neuron[27].syn.SPIKE = {{0, 2}, {0, 3}, {0, 5}, {0, 11}, {0, 12}, {0, 16}, {0, 17}, {0, 20}, {0, 21}, {0, 23}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 31}};
defparam block[0].nb.neuron[28].syn.SPIKE = {{0, 2}, {0, 3}, {0, 4}, {0, 6}, {0, 7}, {0, 9}, {0, 10}, {0, 13}, {0, 14}, {0, 15}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 24}, {0, 25}, {0, 26}, {0, 27}, {0, 29}, {0, 30}};
defparam block[0].nb.neuron[29].syn.SPIKE = {{0, 1}, {0, 4}, {0, 7}, {0, 9}, {0, 10}, {0, 11}, {0, 12}, {0, 13}, {0, 14}, {0, 18}, {0, 19}, {0, 20}, {0, 21}, {0, 22}, {0, 25}, {0, 28}, {0, 30}, {0, 31}};
defparam block[0].nb.neuron[30].syn.SPIKE = {{0, 2}, {0, 3}, {0, 5}, {0, 6}, {0, 10}, {0, 12}, {0, 14}, {0, 15}, {0, 16}, {0, 18}, {0, 19}, {0, 20}, {0, 22}, {0, 23}, {0, 24}, {0, 25}, {0, 26}, {0, 28}, {0, 29}};
defparam block[0].nb.neuron[31].syn.SPIKE = {{0, 1}, {0, 2}, {0, 3}, {0, 4}, {0, 6}, {0, 8}, {0, 9}, {0, 10}, {0, 12}, {0, 14}, {0, 15}, {0, 16}, {0, 17}, {0, 18}, {0, 19}, {0, 22}, {0, 23}, {0, 25}, {0, 27}, {0, 29}};
