// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

interface synapse_if #(WEIGHT=1)
( input clk
, input reset
);
  // --------------------------------------------------------------------
  wire spike;

// --------------------------------------------------------------------
endinterface
