// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

package snn_pkg;

  // --------------------------------------------------------------------
  localparam N = 3; // neurons per block
  localparam T = 2; // number of blocks

  // --------------------------------------------------------------------
  typedef struct {
    int V_0=14;
    int V_REST=6;
    int V_LEAK=1;
    int K_SYN=1;
  } neuron_config_t;

// --------------------------------------------------------------------
endpackage

